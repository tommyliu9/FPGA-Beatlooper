module sinLUT(amount, sinval);
  input [9:0] amount;
  output reg [23:0] sinval;

 always @(amount) begin
   case (amount)
    0: sinval <= 0;
    1: sinval <= 61419;
    2: sinval <= 122835;
    3: sinval <= 184247;
    4: sinval <= 245652;
    5: sinval <= 307048;
    6: sinval <= 368432;
    7: sinval <= 429802;
    8: sinval <= 491156;
    9: sinval <= 552491;
    10: sinval <= 613806;
    11: sinval <= 675097;
    12: sinval <= 736363;
    13: sinval <= 797602;
    14: sinval <= 858810;
    15: sinval <= 919985;
    16: sinval <= 981126;
    17: sinval <= 1042230;
    18: sinval <= 1103295;
    19: sinval <= 1164318;
    20: sinval <= 1225297;
    21: sinval <= 1286230;
    22: sinval <= 1347115;
    23: sinval <= 1407948;
    24: sinval <= 1468729;
    25: sinval <= 1529454;
    26: sinval <= 1590121;
    27: sinval <= 1650728;
    28: sinval <= 1711274;
    29: sinval <= 1771754;
    30: sinval <= 1832168;
    31: sinval <= 1892512;
    32: sinval <= 1952786;
    33: sinval <= 2012985;
    34: sinval <= 2073109;
    35: sinval <= 2133154;
    36: sinval <= 2193119;
    37: sinval <= 2253001;
    38: sinval <= 2312799;
    39: sinval <= 2372509;
    40: sinval <= 2432129;
    41: sinval <= 2491658;
    42: sinval <= 2551092;
    43: sinval <= 2610431;
    44: sinval <= 2669671;
    45: sinval <= 2728810;
    46: sinval <= 2787847;
    47: sinval <= 2846778;
    48: sinval <= 2905602;
    49: sinval <= 2964316;
    50: sinval <= 3022918;
    51: sinval <= 3081407;
    52: sinval <= 3139779;
    53: sinval <= 3198032;
    54: sinval <= 3256165;
    55: sinval <= 3314176;
    56: sinval <= 3372061;
    57: sinval <= 3429819;
    58: sinval <= 3487447;
    59: sinval <= 3544944;
    60: sinval <= 3602308;
    61: sinval <= 3659535;
    62: sinval <= 3716625;
    63: sinval <= 3773574;
    64: sinval <= 3830381;
    65: sinval <= 3887043;
    66: sinval <= 3943559;
    67: sinval <= 3999925;
    68: sinval <= 4056142;
    69: sinval <= 4112205;
    70: sinval <= 4168112;
    71: sinval <= 4223863;
    72: sinval <= 4279454;
    73: sinval <= 4334884;
    74: sinval <= 4390151;
    75: sinval <= 4445251;
    76: sinval <= 4500185;
    77: sinval <= 4554948;
    78: sinval <= 4609539;
    79: sinval <= 4663957;
    80: sinval <= 4718199;
    81: sinval <= 4772262;
    82: sinval <= 4826146;
    83: sinval <= 4879848;
    84: sinval <= 4933365;
    85: sinval <= 4986696;
    86: sinval <= 5039840;
    87: sinval <= 5092793;
    88: sinval <= 5145554;
    89: sinval <= 5198121;
    90: sinval <= 5250492;
    91: sinval <= 5302665;
    92: sinval <= 5354637;
    93: sinval <= 5406408;
    94: sinval <= 5457975;
    95: sinval <= 5509336;
    96: sinval <= 5560489;
    97: sinval <= 5611432;
    98: sinval <= 5662164;
    99: sinval <= 5712682;
    100: sinval <= 5762985;
    101: sinval <= 5813070;
    102: sinval <= 5862936;
    103: sinval <= 5912581;
    104: sinval <= 5962002;
    105: sinval <= 6011199;
    106: sinval <= 6060169;
    107: sinval <= 6108910;
    108: sinval <= 6157421;
    109: sinval <= 6205700;
    110: sinval <= 6253745;
    111: sinval <= 6301553;
    112: sinval <= 6349124;
    113: sinval <= 6396456;
    114: sinval <= 6443546;
    115: sinval <= 6490393;
    116: sinval <= 6536995;
    117: sinval <= 6583351;
    118: sinval <= 6629458;
    119: sinval <= 6675315;
    120: sinval <= 6720921;
    121: sinval <= 6766273;
    122: sinval <= 6811369;
    123: sinval <= 6856209;
    124: sinval <= 6900790;
    125: sinval <= 6945111;
    126: sinval <= 6989170;
    127: sinval <= 7032965;
    128: sinval <= 7076494;
    129: sinval <= 7119757;
    130: sinval <= 7162752;
    131: sinval <= 7205476;
    132: sinval <= 7247928;
    133: sinval <= 7290107;
    134: sinval <= 7332011;
    135: sinval <= 7373638;
    136: sinval <= 7414987;
    137: sinval <= 7456056;
    138: sinval <= 7496844;
    139: sinval <= 7537350;
    140: sinval <= 7577571;
    141: sinval <= 7617506;
    142: sinval <= 7657153;
    143: sinval <= 7696512;
    144: sinval <= 7735581;
    145: sinval <= 7774358;
    146: sinval <= 7812841;
    147: sinval <= 7851030;
    148: sinval <= 7888923;
    149: sinval <= 7926518;
    150: sinval <= 7963814;
    151: sinval <= 8000809;
    152: sinval <= 8037503;
    153: sinval <= 8073893;
    154: sinval <= 8109979;
    155: sinval <= 8145760;
    156: sinval <= 8181232;
    157: sinval <= 8216396;
    158: sinval <= 8251251;
    159: sinval <= 8285794;
    160: sinval <= 8320024;
    161: sinval <= 8353940;
    162: sinval <= 8387542;
    163: sinval <= 8420827;
    164: sinval <= 8453794;
    165: sinval <= 8486443;
    166: sinval <= 8518771;
    167: sinval <= 8550778;
    168: sinval <= 8582462;
    169: sinval <= 8613823;
    170: sinval <= 8644858;
    171: sinval <= 8675568;
    172: sinval <= 8705950;
    173: sinval <= 8736004;
    174: sinval <= 8765728;
    175: sinval <= 8795122;
    176: sinval <= 8824184;
    177: sinval <= 8852913;
    178: sinval <= 8881308;
    179: sinval <= 8909368;
    180: sinval <= 8937092;
    181: sinval <= 8964479;
    182: sinval <= 8991527;
    183: sinval <= 9018237;
    184: sinval <= 9044606;
    185: sinval <= 9070634;
    186: sinval <= 9096320;
    187: sinval <= 9121663;
    188: sinval <= 9146661;
    189: sinval <= 9171315;
    190: sinval <= 9195623;
    191: sinval <= 9219583;
    192: sinval <= 9243196;
    193: sinval <= 9266460;
    194: sinval <= 9289375;
    195: sinval <= 9311939;
    196: sinval <= 9334152;
    197: sinval <= 9356013;
    198: sinval <= 9377521;
    199: sinval <= 9398676;
    200: sinval <= 9419475;
    201: sinval <= 9439920;
    202: sinval <= 9460008;
    203: sinval <= 9479739;
    204: sinval <= 9499113;
    205: sinval <= 9518128;
    206: sinval <= 9536785;
    207: sinval <= 9555081;
    208: sinval <= 9573017;
    209: sinval <= 9590592;
    210: sinval <= 9607806;
    211: sinval <= 9624657;
    212: sinval <= 9641144;
    213: sinval <= 9657268;
    214: sinval <= 9673028;
    215: sinval <= 9688423;
    216: sinval <= 9703452;
    217: sinval <= 9718116;
    218: sinval <= 9732412;
    219: sinval <= 9746342;
    220: sinval <= 9759904;
    221: sinval <= 9773098;
    222: sinval <= 9785923;
    223: sinval <= 9798379;
    224: sinval <= 9810465;
    225: sinval <= 9822181;
    226: sinval <= 9833527;
    227: sinval <= 9844502;
    228: sinval <= 9855105;
    229: sinval <= 9865337;
    230: sinval <= 9875196;
    231: sinval <= 9884683;
    232: sinval <= 9893797;
    233: sinval <= 9902538;
    234: sinval <= 9910905;
    235: sinval <= 9918899;
    236: sinval <= 9926518;
    237: sinval <= 9933763;
    238: sinval <= 9940633;
    239: sinval <= 9947128;
    240: sinval <= 9953248;
    241: sinval <= 9958992;
    242: sinval <= 9964361;
    243: sinval <= 9969354;
    244: sinval <= 9973971;
    245: sinval <= 9978211;
    246: sinval <= 9982075;
    247: sinval <= 9985563;
    248: sinval <= 9988673;
    249: sinval <= 9991407;
    250: sinval <= 9993765;
    251: sinval <= 9995745;
    252: sinval <= 9997348;
    253: sinval <= 9998574;
    254: sinval <= 9999422;
    255: sinval <= 9999894;
    256: sinval <= 9999988;
    257: sinval <= 9999705;
    258: sinval <= 9999045;
    259: sinval <= 9998008;
    260: sinval <= 9996593;
    261: sinval <= 9994802;
    262: sinval <= 9992633;
    263: sinval <= 9990088;
    264: sinval <= 9987165;
    265: sinval <= 9983866;
    266: sinval <= 9980190;
    267: sinval <= 9976138;
    268: sinval <= 9971709;
    269: sinval <= 9966904;
    270: sinval <= 9961724;
    271: sinval <= 9956167;
    272: sinval <= 9950235;
    273: sinval <= 9943927;
    274: sinval <= 9937245;
    275: sinval <= 9930187;
    276: sinval <= 9922755;
    277: sinval <= 9914949;
    278: sinval <= 9906769;
    279: sinval <= 9898214;
    280: sinval <= 9889287;
    281: sinval <= 9879986;
    282: sinval <= 9870313;
    283: sinval <= 9860267;
    284: sinval <= 9849850;
    285: sinval <= 9839061;
    286: sinval <= 9827901;
    287: sinval <= 9816369;
    288: sinval <= 9804468;
    289: sinval <= 9792197;
    290: sinval <= 9779556;
    291: sinval <= 9766547;
    292: sinval <= 9753169;
    293: sinval <= 9739423;
    294: sinval <= 9725310;
    295: sinval <= 9710830;
    296: sinval <= 9695983;
    297: sinval <= 9680771;
    298: sinval <= 9665194;
    299: sinval <= 9649252;
    300: sinval <= 9632946;
    301: sinval <= 9616276;
    302: sinval <= 9599244;
    303: sinval <= 9581850;
    304: sinval <= 9564094;
    305: sinval <= 9545978;
    306: sinval <= 9527501;
    307: sinval <= 9508665;
    308: sinval <= 9489471;
    309: sinval <= 9469918;
    310: sinval <= 9450008;
    311: sinval <= 9429742;
    312: sinval <= 9409120;
    313: sinval <= 9388143;
    314: sinval <= 9366812;
    315: sinval <= 9345127;
    316: sinval <= 9323090;
    317: sinval <= 9300701;
    318: sinval <= 9277962;
    319: sinval <= 9254872;
    320: sinval <= 9231433;
    321: sinval <= 9207646;
    322: sinval <= 9183512;
    323: sinval <= 9159031;
    324: sinval <= 9134205;
    325: sinval <= 9109034;
    326: sinval <= 9083520;
    327: sinval <= 9057663;
    328: sinval <= 9031464;
    329: sinval <= 9004925;
    330: sinval <= 8978045;
    331: sinval <= 8950828;
    332: sinval <= 8923272;
    333: sinval <= 8895380;
    334: sinval <= 8867152;
    335: sinval <= 8838590;
    336: sinval <= 8809695;
    337: sinval <= 8780467;
    338: sinval <= 8750908;
    339: sinval <= 8721018;
    340: sinval <= 8690800;
    341: sinval <= 8660254;
    342: sinval <= 8629381;
    343: sinval <= 8598183;
    344: sinval <= 8566660;
    345: sinval <= 8534815;
    346: sinval <= 8502647;
    347: sinval <= 8470158;
    348: sinval <= 8437350;
    349: sinval <= 8404224;
    350: sinval <= 8370781;
    351: sinval <= 8337022;
    352: sinval <= 8302948;
    353: sinval <= 8268561;
    354: sinval <= 8233862;
    355: sinval <= 8198853;
    356: sinval <= 8163534;
    357: sinval <= 8127908;
    358: sinval <= 8091975;
    359: sinval <= 8055736;
    360: sinval <= 8019194;
    361: sinval <= 7982349;
    362: sinval <= 7945203;
    363: sinval <= 7907757;
    364: sinval <= 7870013;
    365: sinval <= 7831973;
    366: sinval <= 7793636;
    367: sinval <= 7755006;
    368: sinval <= 7716083;
    369: sinval <= 7676869;
    370: sinval <= 7637366;
    371: sinval <= 7597574;
    372: sinval <= 7557496;
    373: sinval <= 7517132;
    374: sinval <= 7476486;
    375: sinval <= 7435557;
    376: sinval <= 7394347;
    377: sinval <= 7352859;
    378: sinval <= 7311093;
    379: sinval <= 7269052;
    380: sinval <= 7226736;
    381: sinval <= 7184147;
    382: sinval <= 7141288;
    383: sinval <= 7098159;
    384: sinval <= 7054763;
    385: sinval <= 7011100;
    386: sinval <= 6967173;
    387: sinval <= 6922983;
    388: sinval <= 6878532;
    389: sinval <= 6833821;
    390: sinval <= 6788853;
    391: sinval <= 6743629;
    392: sinval <= 6698150;
    393: sinval <= 6652418;
    394: sinval <= 6606436;
    395: sinval <= 6560204;
    396: sinval <= 6513725;
    397: sinval <= 6467000;
    398: sinval <= 6420031;
    399: sinval <= 6372820;
    400: sinval <= 6325369;
    401: sinval <= 6277679;
    402: sinval <= 6229752;
    403: sinval <= 6181590;
    404: sinval <= 6133195;
    405: sinval <= 6084568;
    406: sinval <= 6035712;
    407: sinval <= 5986629;
    408: sinval <= 5937319;
    409: sinval <= 5887786;
    410: sinval <= 5838030;
    411: sinval <= 5788055;
    412: sinval <= 5737860;
    413: sinval <= 5687450;
    414: sinval <= 5636825;
    415: sinval <= 5585987;
    416: sinval <= 5534939;
    417: sinval <= 5483681;
    418: sinval <= 5432217;
    419: sinval <= 5380548;
    420: sinval <= 5328676;
    421: sinval <= 5276603;
    422: sinval <= 5224331;
    423: sinval <= 5171862;
    424: sinval <= 5119198;
    425: sinval <= 5066340;
    426: sinval <= 5013292;
    427: sinval <= 4960054;
    428: sinval <= 4906629;
    429: sinval <= 4853020;
    430: sinval <= 4799227;
    431: sinval <= 4745253;
    432: sinval <= 4691100;
    433: sinval <= 4636770;
    434: sinval <= 4582265;
    435: sinval <= 4527588;
    436: sinval <= 4472739;
    437: sinval <= 4417722;
    438: sinval <= 4362538;
    439: sinval <= 4307190;
    440: sinval <= 4251679;
    441: sinval <= 4196008;
    442: sinval <= 4140178;
    443: sinval <= 4084192;
    444: sinval <= 4028052;
    445: sinval <= 3971761;
    446: sinval <= 3915319;
    447: sinval <= 3858730;
    448: sinval <= 3801995;
    449: sinval <= 3745117;
    450: sinval <= 3688097;
    451: sinval <= 3630939;
    452: sinval <= 3573643;
    453: sinval <= 3516213;
    454: sinval <= 3458649;
    455: sinval <= 3400956;
    456: sinval <= 3343134;
    457: sinval <= 3285186;
    458: sinval <= 3227114;
    459: sinval <= 3168921;
    460: sinval <= 3110607;
    461: sinval <= 3052177;
    462: sinval <= 2993631;
    463: sinval <= 2934973;
    464: sinval <= 2876203;
    465: sinval <= 2817326;
    466: sinval <= 2758341;
    467: sinval <= 2699253;
    468: sinval <= 2640063;
    469: sinval <= 2580774;
    470: sinval <= 2521387;
    471: sinval <= 2461905;
    472: sinval <= 2402330;
    473: sinval <= 2342665;
    474: sinval <= 2282911;
    475: sinval <= 2223071;
    476: sinval <= 2163147;
    477: sinval <= 2103141;
    478: sinval <= 2043057;
    479: sinval <= 1982895;
    480: sinval <= 1922658;
    481: sinval <= 1862349;
    482: sinval <= 1801969;
    483: sinval <= 1741522;
    484: sinval <= 1681009;
    485: sinval <= 1620432;
    486: sinval <= 1559795;
    487: sinval <= 1499098;
    488: sinval <= 1438345;
    489: sinval <= 1377538;
    490: sinval <= 1316679;
    491: sinval <= 1255770;
    492: sinval <= 1194813;
    493: sinval <= 1133812;
    494: sinval <= 1072768;
    495: sinval <= 1011683;
    496: sinval <= 950560;
    497: sinval <= 889402;
    498: sinval <= 828210;
    499: sinval <= 766986;
    500: sinval <= 705734;
    501: sinval <= 644455;
    502: sinval <= 583151;
    503: sinval <= 521826;
    504: sinval <= 460481;
    505: sinval <= 399119;
    506: sinval <= 337741;
    507: sinval <= 276351;
    508: sinval <= 214951;
    509: sinval <= 153542;
    510: sinval <= 92128;
    511: sinval <= 30710;
    512: sinval <= -30710;
    513: sinval <= -92128;
    514: sinval <= -153542;
    515: sinval <= -214951;
    516: sinval <= -276351;
    517: sinval <= -337741;
    518: sinval <= -399119;
    519: sinval <= -460481;
    520: sinval <= -521826;
    521: sinval <= -583151;
    522: sinval <= -644455;
    523: sinval <= -705734;
    524: sinval <= -766986;
    525: sinval <= -828210;
    526: sinval <= -889402;
    527: sinval <= -950560;
    528: sinval <= -1011683;
    529: sinval <= -1072768;
    530: sinval <= -1133812;
    531: sinval <= -1194813;
    532: sinval <= -1255770;
    533: sinval <= -1316679;
    534: sinval <= -1377538;
    535: sinval <= -1438345;
    536: sinval <= -1499098;
    537: sinval <= -1559795;
    538: sinval <= -1620432;
    539: sinval <= -1681009;
    540: sinval <= -1741522;
    541: sinval <= -1801969;
    542: sinval <= -1862349;
    543: sinval <= -1922658;
    544: sinval <= -1982895;
    545: sinval <= -2043057;
    546: sinval <= -2103141;
    547: sinval <= -2163147;
    548: sinval <= -2223071;
    549: sinval <= -2282911;
    550: sinval <= -2342665;
    551: sinval <= -2402330;
    552: sinval <= -2461905;
    553: sinval <= -2521387;
    554: sinval <= -2580774;
    555: sinval <= -2640063;
    556: sinval <= -2699253;
    557: sinval <= -2758341;
    558: sinval <= -2817326;
    559: sinval <= -2876203;
    560: sinval <= -2934973;
    561: sinval <= -2993631;
    562: sinval <= -3052177;
    563: sinval <= -3110607;
    564: sinval <= -3168921;
    565: sinval <= -3227114;
    566: sinval <= -3285186;
    567: sinval <= -3343134;
    568: sinval <= -3400956;
    569: sinval <= -3458649;
    570: sinval <= -3516213;
    571: sinval <= -3573643;
    572: sinval <= -3630939;
    573: sinval <= -3688097;
    574: sinval <= -3745117;
    575: sinval <= -3801995;
    576: sinval <= -3858730;
    577: sinval <= -3915319;
    578: sinval <= -3971761;
    579: sinval <= -4028052;
    580: sinval <= -4084192;
    581: sinval <= -4140178;
    582: sinval <= -4196008;
    583: sinval <= -4251679;
    584: sinval <= -4307190;
    585: sinval <= -4362538;
    586: sinval <= -4417722;
    587: sinval <= -4472739;
    588: sinval <= -4527588;
    589: sinval <= -4582265;
    590: sinval <= -4636770;
    591: sinval <= -4691100;
    592: sinval <= -4745253;
    593: sinval <= -4799227;
    594: sinval <= -4853020;
    595: sinval <= -4906629;
    596: sinval <= -4960054;
    597: sinval <= -5013292;
    598: sinval <= -5066340;
    599: sinval <= -5119198;
    600: sinval <= -5171862;
    601: sinval <= -5224331;
    602: sinval <= -5276603;
    603: sinval <= -5328676;
    604: sinval <= -5380548;
    605: sinval <= -5432217;
    606: sinval <= -5483681;
    607: sinval <= -5534939;
    608: sinval <= -5585987;
    609: sinval <= -5636825;
    610: sinval <= -5687450;
    611: sinval <= -5737860;
    612: sinval <= -5788055;
    613: sinval <= -5838030;
    614: sinval <= -5887786;
    615: sinval <= -5937319;
    616: sinval <= -5986629;
    617: sinval <= -6035712;
    618: sinval <= -6084568;
    619: sinval <= -6133195;
    620: sinval <= -6181590;
    621: sinval <= -6229752;
    622: sinval <= -6277679;
    623: sinval <= -6325369;
    624: sinval <= -6372820;
    625: sinval <= -6420031;
    626: sinval <= -6467000;
    627: sinval <= -6513725;
    628: sinval <= -6560204;
    629: sinval <= -6606436;
    630: sinval <= -6652418;
    631: sinval <= -6698150;
    632: sinval <= -6743629;
    633: sinval <= -6788853;
    634: sinval <= -6833821;
    635: sinval <= -6878532;
    636: sinval <= -6922983;
    637: sinval <= -6967173;
    638: sinval <= -7011100;
    639: sinval <= -7054763;
    640: sinval <= -7098159;
    641: sinval <= -7141288;
    642: sinval <= -7184147;
    643: sinval <= -7226736;
    644: sinval <= -7269052;
    645: sinval <= -7311093;
    646: sinval <= -7352859;
    647: sinval <= -7394347;
    648: sinval <= -7435557;
    649: sinval <= -7476486;
    650: sinval <= -7517132;
    651: sinval <= -7557496;
    652: sinval <= -7597574;
    653: sinval <= -7637366;
    654: sinval <= -7676869;
    655: sinval <= -7716083;
    656: sinval <= -7755006;
    657: sinval <= -7793636;
    658: sinval <= -7831973;
    659: sinval <= -7870013;
    660: sinval <= -7907757;
    661: sinval <= -7945203;
    662: sinval <= -7982349;
    663: sinval <= -8019194;
    664: sinval <= -8055736;
    665: sinval <= -8091975;
    666: sinval <= -8127908;
    667: sinval <= -8163534;
    668: sinval <= -8198853;
    669: sinval <= -8233862;
    670: sinval <= -8268561;
    671: sinval <= -8302948;
    672: sinval <= -8337022;
    673: sinval <= -8370781;
    674: sinval <= -8404224;
    675: sinval <= -8437350;
    676: sinval <= -8470158;
    677: sinval <= -8502647;
    678: sinval <= -8534815;
    679: sinval <= -8566660;
    680: sinval <= -8598183;
    681: sinval <= -8629381;
    682: sinval <= -8660254;
    683: sinval <= -8690800;
    684: sinval <= -8721018;
    685: sinval <= -8750908;
    686: sinval <= -8780467;
    687: sinval <= -8809695;
    688: sinval <= -8838590;
    689: sinval <= -8867152;
    690: sinval <= -8895380;
    691: sinval <= -8923272;
    692: sinval <= -8950828;
    693: sinval <= -8978045;
    694: sinval <= -9004925;
    695: sinval <= -9031464;
    696: sinval <= -9057663;
    697: sinval <= -9083520;
    698: sinval <= -9109034;
    699: sinval <= -9134205;
    700: sinval <= -9159031;
    701: sinval <= -9183512;
    702: sinval <= -9207646;
    703: sinval <= -9231433;
    704: sinval <= -9254872;
    705: sinval <= -9277962;
    706: sinval <= -9300701;
    707: sinval <= -9323090;
    708: sinval <= -9345127;
    709: sinval <= -9366812;
    710: sinval <= -9388143;
    711: sinval <= -9409120;
    712: sinval <= -9429742;
    713: sinval <= -9450008;
    714: sinval <= -9469918;
    715: sinval <= -9489471;
    716: sinval <= -9508665;
    717: sinval <= -9527501;
    718: sinval <= -9545978;
    719: sinval <= -9564094;
    720: sinval <= -9581850;
    721: sinval <= -9599244;
    722: sinval <= -9616276;
    723: sinval <= -9632946;
    724: sinval <= -9649252;
    725: sinval <= -9665194;
    726: sinval <= -9680771;
    727: sinval <= -9695983;
    728: sinval <= -9710830;
    729: sinval <= -9725310;
    730: sinval <= -9739423;
    731: sinval <= -9753169;
    732: sinval <= -9766547;
    733: sinval <= -9779556;
    734: sinval <= -9792197;
    735: sinval <= -9804468;
    736: sinval <= -9816369;
    737: sinval <= -9827901;
    738: sinval <= -9839061;
    739: sinval <= -9849850;
    740: sinval <= -9860267;
    741: sinval <= -9870313;
    742: sinval <= -9879986;
    743: sinval <= -9889287;
    744: sinval <= -9898214;
    745: sinval <= -9906769;
    746: sinval <= -9914949;
    747: sinval <= -9922755;
    748: sinval <= -9930187;
    749: sinval <= -9937245;
    750: sinval <= -9943927;
    751: sinval <= -9950235;
    752: sinval <= -9956167;
    753: sinval <= -9961724;
    754: sinval <= -9966904;
    755: sinval <= -9971709;
    756: sinval <= -9976138;
    757: sinval <= -9980190;
    758: sinval <= -9983866;
    759: sinval <= -9987165;
    760: sinval <= -9990088;
    761: sinval <= -9992633;
    762: sinval <= -9994802;
    763: sinval <= -9996593;
    764: sinval <= -9998008;
    765: sinval <= -9999045;
    766: sinval <= -9999705;
    767: sinval <= -9999988;
    768: sinval <= -9999894;
    769: sinval <= -9999422;
    770: sinval <= -9998574;
    771: sinval <= -9997348;
    772: sinval <= -9995745;
    773: sinval <= -9993765;
    774: sinval <= -9991407;
    775: sinval <= -9988673;
    776: sinval <= -9985563;
    777: sinval <= -9982075;
    778: sinval <= -9978211;
    779: sinval <= -9973971;
    780: sinval <= -9969354;
    781: sinval <= -9964361;
    782: sinval <= -9958992;
    783: sinval <= -9953248;
    784: sinval <= -9947128;
    785: sinval <= -9940633;
    786: sinval <= -9933763;
    787: sinval <= -9926518;
    788: sinval <= -9918899;
    789: sinval <= -9910905;
    790: sinval <= -9902538;
    791: sinval <= -9893797;
    792: sinval <= -9884683;
    793: sinval <= -9875196;
    794: sinval <= -9865337;
    795: sinval <= -9855105;
    796: sinval <= -9844502;
    797: sinval <= -9833527;
    798: sinval <= -9822181;
    799: sinval <= -9810465;
    800: sinval <= -9798379;
    801: sinval <= -9785923;
    802: sinval <= -9773098;
    803: sinval <= -9759904;
    804: sinval <= -9746342;
    805: sinval <= -9732412;
    806: sinval <= -9718116;
    807: sinval <= -9703452;
    808: sinval <= -9688423;
    809: sinval <= -9673028;
    810: sinval <= -9657268;
    811: sinval <= -9641144;
    812: sinval <= -9624657;
    813: sinval <= -9607806;
    814: sinval <= -9590592;
    815: sinval <= -9573017;
    816: sinval <= -9555081;
    817: sinval <= -9536785;
    818: sinval <= -9518128;
    819: sinval <= -9499113;
    820: sinval <= -9479739;
    821: sinval <= -9460008;
    822: sinval <= -9439920;
    823: sinval <= -9419475;
    824: sinval <= -9398676;
    825: sinval <= -9377521;
    826: sinval <= -9356013;
    827: sinval <= -9334152;
    828: sinval <= -9311939;
    829: sinval <= -9289375;
    830: sinval <= -9266460;
    831: sinval <= -9243196;
    832: sinval <= -9219583;
    833: sinval <= -9195623;
    834: sinval <= -9171315;
    835: sinval <= -9146661;
    836: sinval <= -9121663;
    837: sinval <= -9096320;
    838: sinval <= -9070634;
    839: sinval <= -9044606;
    840: sinval <= -9018237;
    841: sinval <= -8991527;
    842: sinval <= -8964479;
    843: sinval <= -8937092;
    844: sinval <= -8909368;
    845: sinval <= -8881308;
    846: sinval <= -8852913;
    847: sinval <= -8824184;
    848: sinval <= -8795122;
    849: sinval <= -8765728;
    850: sinval <= -8736004;
    851: sinval <= -8705950;
    852: sinval <= -8675568;
    853: sinval <= -8644858;
    854: sinval <= -8613823;
    855: sinval <= -8582462;
    856: sinval <= -8550778;
    857: sinval <= -8518771;
    858: sinval <= -8486443;
    859: sinval <= -8453794;
    860: sinval <= -8420827;
    861: sinval <= -8387542;
    862: sinval <= -8353940;
    863: sinval <= -8320024;
    864: sinval <= -8285794;
    865: sinval <= -8251251;
    866: sinval <= -8216396;
    867: sinval <= -8181232;
    868: sinval <= -8145760;
    869: sinval <= -8109979;
    870: sinval <= -8073893;
    871: sinval <= -8037503;
    872: sinval <= -8000809;
    873: sinval <= -7963814;
    874: sinval <= -7926518;
    875: sinval <= -7888923;
    876: sinval <= -7851030;
    877: sinval <= -7812841;
    878: sinval <= -7774358;
    879: sinval <= -7735581;
    880: sinval <= -7696512;
    881: sinval <= -7657153;
    882: sinval <= -7617506;
    883: sinval <= -7577571;
    884: sinval <= -7537350;
    885: sinval <= -7496844;
    886: sinval <= -7456056;
    887: sinval <= -7414987;
    888: sinval <= -7373638;
    889: sinval <= -7332011;
    890: sinval <= -7290107;
    891: sinval <= -7247928;
    892: sinval <= -7205476;
    893: sinval <= -7162752;
    894: sinval <= -7119757;
    895: sinval <= -7076494;
    896: sinval <= -7032965;
    897: sinval <= -6989170;
    898: sinval <= -6945111;
    899: sinval <= -6900790;
    900: sinval <= -6856209;
    901: sinval <= -6811369;
    902: sinval <= -6766273;
    903: sinval <= -6720921;
    904: sinval <= -6675315;
    905: sinval <= -6629458;
    906: sinval <= -6583351;
    907: sinval <= -6536995;
    908: sinval <= -6490393;
    909: sinval <= -6443546;
    910: sinval <= -6396456;
    911: sinval <= -6349124;
    912: sinval <= -6301553;
    913: sinval <= -6253745;
    914: sinval <= -6205700;
    915: sinval <= -6157421;
    916: sinval <= -6108910;
    917: sinval <= -6060169;
    918: sinval <= -6011199;
    919: sinval <= -5962002;
    920: sinval <= -5912581;
    921: sinval <= -5862936;
    922: sinval <= -5813070;
    923: sinval <= -5762985;
    924: sinval <= -5712682;
    925: sinval <= -5662164;
    926: sinval <= -5611432;
    927: sinval <= -5560489;
    928: sinval <= -5509336;
    929: sinval <= -5457975;
    930: sinval <= -5406408;
    931: sinval <= -5354637;
    932: sinval <= -5302665;
    933: sinval <= -5250492;
    934: sinval <= -5198121;
    935: sinval <= -5145554;
    936: sinval <= -5092793;
    937: sinval <= -5039840;
    938: sinval <= -4986696;
    939: sinval <= -4933365;
    940: sinval <= -4879848;
    941: sinval <= -4826146;
    942: sinval <= -4772262;
    943: sinval <= -4718199;
    944: sinval <= -4663957;
    945: sinval <= -4609539;
    946: sinval <= -4554948;
    947: sinval <= -4500185;
    948: sinval <= -4445251;
    949: sinval <= -4390151;
    950: sinval <= -4334884;
    951: sinval <= -4279454;
    952: sinval <= -4223863;
    953: sinval <= -4168112;
    954: sinval <= -4112205;
    955: sinval <= -4056142;
    956: sinval <= -3999925;
    957: sinval <= -3943559;
    958: sinval <= -3887043;
    959: sinval <= -3830381;
    960: sinval <= -3773574;
    961: sinval <= -3716625;
    962: sinval <= -3659535;
    963: sinval <= -3602308;
    964: sinval <= -3544944;
    965: sinval <= -3487447;
    966: sinval <= -3429819;
    967: sinval <= -3372061;
    968: sinval <= -3314176;
    969: sinval <= -3256165;
    970: sinval <= -3198032;
    971: sinval <= -3139779;
    972: sinval <= -3081407;
    973: sinval <= -3022918;
    974: sinval <= -2964316;
    975: sinval <= -2905602;
    976: sinval <= -2846778;
    977: sinval <= -2787847;
    978: sinval <= -2728810;
    979: sinval <= -2669671;
    980: sinval <= -2610431;
    981: sinval <= -2551092;
    982: sinval <= -2491658;
    983: sinval <= -2432129;
    984: sinval <= -2372509;
    985: sinval <= -2312799;
    986: sinval <= -2253001;
    987: sinval <= -2193119;
    988: sinval <= -2133154;
    989: sinval <= -2073109;
    990: sinval <= -2012985;
    991: sinval <= -1952786;
    992: sinval <= -1892512;
    993: sinval <= -1832168;
    994: sinval <= -1771754;
    995: sinval <= -1711274;
    996: sinval <= -1650728;
    997: sinval <= -1590121;
    998: sinval <= -1529454;
    999: sinval <= -1468729;
    1000: sinval <= -1407948;
    1001: sinval <= -1347115;
    1002: sinval <= -1286230;
    1003: sinval <= -1225297;
    1004: sinval <= -1164318;
    1005: sinval <= -1103295;
    1006: sinval <= -1042230;
    1007: sinval <= -981126;
    1008: sinval <= -919985;
    1009: sinval <= -858810;
    1010: sinval <= -797602;
    1011: sinval <= -736363;
    1012: sinval <= -675097;
    1013: sinval <= -613806;
    1014: sinval <= -552491;
    1015: sinval <= -491156;
    1016: sinval <= -429802;
    1017: sinval <= -368432;
    1018: sinval <= -307048;
    1019: sinval <= -245652;
    1020: sinval <= -184247;
    1021: sinval <= -122835;
    1022: sinval <= -61419;
    1023: sinval <= 0;
	 default: sinval <= 0;
   endcase
  end

endmodule
